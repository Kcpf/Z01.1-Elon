-- Elementos de Sistemas
-- by Luciano Soares
-- HalfAdder.vhd

-- Implementa Half Adder

Library ieee;
use ieee.std_logic_1164.all;

entity HalfAdder is
	port(
		a,b:         in STD_LOGIC;   -- entradas
		soma,vaium: out STD_LOGIC   -- sum e carry
	);
end entity;

architecture rtl of HalfAdder is
  -- Aqui declaramos sinais (fios auxiliares)
  -- e componentes (outros módulos) que serao
  -- utilizados nesse modulo.

begin
<<<<<<< HEAD
  soma <= a xor b;
  vaium <= a and b;
=======
  -- Implementação vem aqui!
	soma <= a xor b;
	vaium <= a and b;
>>>>>>> 0c675ccf355e2c8c18fe25ee4847eb1a921fd42c

end architecture;
