-- Elementos de Sistemas
-- developed by Luciano Soares
-- file: tb_ALU.vhd
-- date: 4/4/2017

library ieee;
use ieee.std_logic_1164.all;

library vunit_lib;
context vunit_lib.vunit_context;

entity tb_ALU is
  generic (runner_cfg : string);
end entity;

architecture tb of tb_ALU is

component ALU is
	port (
    x,y:   in STD_LOGIC_VECTOR(15 downto 0); -- entradas de dados da ALU
    zx:    in STD_LOGIC;                     -- zera a entrada x
    nx:    in STD_LOGIC;                     -- inverte a entrada x
    sizex: in STD_LOGIC_VECTOR(2 downto 0);  -- tamanho do shift em x
    dirx:  in STD_LOGIC;                     -- direcao do shift em x
    zy:    in STD_LOGIC;                     -- zera a entrada y
    ny:    in STD_LOGIC;                     -- inverte a entrada y
    sizey: in STD_LOGIC_VECTOR(2 downto 0);  -- tamanho do shift em y
    diry:  in STD_LOGIC;                     -- direcao do shift em y
    f:     in STD_LOGIC_VECTOR(1 downto 0);  -- se 0 calcula x & y, senão x + y
    no:    in STD_LOGIC;                     -- inverte o valor da saída
    zr:    out STD_LOGIC;                    -- setado se saída igual a zero
    ng:    out STD_LOGIC;                    -- setado se saída é negativa
    carry: out STD_LOGIC;                    -- carry da soma
    saida: out STD_LOGIC_VECTOR(15 downto 0) -- saída de dados da ALU
	);
end component;

   signal  inX, inY : STD_LOGIC_VECTOR(15 downto 0);
   signal  inF : STD_LOGIC_VECTOR(1 downto 0);
   signal  inSizeX, inSizeY : STD_LOGIC_VECTOR(2 downto 0);
   signal  inZX, inNX, inZY, inNY, inNO, outZR, outNG, outCA, inDirX, inDirY : STD_LOGIC;
   signal  outSaida : STD_LOGIC_VECTOR(15 downto 0);

begin

	mapping: ALU port map(
    x  => inX,
    y  => inY,
    zx => inZx,
    nx => inNx,
    sizex => inSizeX,
    dirx => inDirX,
    zy => inZy,
    ny => inNy,
    sizey => inSizeY,
    diry => inDirY,
    f  => inF,
    no => inNo,
    zr => outZr,
    ng => outNg,
    carry => outCa,
    saida => outsaida);

  main : process
  begin
    test_runner_setup(runner, runner_cfg);

      -- Teste: 1
      inX <= "0000000000000000"; inY <= "1111111111111111";
      inZX <= '1'; inNX <= '0'; inZY <= '1'; inNY <= '0'; inF <= "01"; inNO <= '0'; inSizeX <= "000"; inSizeY <= "000"; inDirX <= '0'; inDirY <= '0';
      wait for 100 ps;
      assert(outZR = '1' and outNG = '0' and outSaida= "0000000000000000")  report "Falha em teste: 1" severity error;

      -- Teste: 2
      inX <= "0000000000000000"; inY <= "1111111111111111";
      inZX <= '1'; inNX <= '1'; inZY <= '1'; inNY <= '1'; inF <= "01"; inNO <= '1'; inSizeX <= "000"; inSizeY <= "000"; inDirX <= '0'; inDirY <= '0';
      wait for 200 ps;
      assert(outZR = '0' and outNG = '0' and outSaida= "0000000000000001")  report "Falha em teste: 2" severity error;

      -- Teste: 3
      inX <= "0000000000000000"; inY <= "1111111111111111";
      inZX <= '1'; inNX <= '1'; inZY <= '1'; inNY <= '0'; inF <= "01"; inNO <= '0'; inSizeX <= "000"; inSizeY <= "000"; inDirX <= '0'; inDirY <= '0';
      wait for 200 ps;
      assert(outZR = '0' and outNG = '1' and outSaida= "1111111111111111")  report "Falha em teste: 3" severity error;

      -- Teste: 4
      inX <= "0000000000000000"; inY <= "1111111111111111";
      inZX <= '0'; inNX <= '0'; inZY <= '1'; inNY <= '1'; inF <= "00"; inNO <= '0'; inSizeX <= "000"; inSizeY <= "000"; inDirX <= '0'; inDirY <= '0';
      wait for 200 ps;
      assert(outZR = '1' and outNG = '0' and outSaida= "0000000000000000")  report "Falha em teste: 4" severity error;

      -- Teste: 5
      inX <= "0000000000000000"; inY <= "1111111111111111";
      inZX <= '1'; inNX <= '1'; inZY <= '0'; inNY <= '0'; inF <= "00"; inNO <= '0'; inSizeX <= "000"; inSizeY <= "000"; inDirX <= '0'; inDirY <= '0';
      wait for 200 ps;
      assert(outZR = '0' and outNG = '1' and outSaida= "1111111111111111")  report "Falha em teste: 5" severity error;

      -- Teste: 6
      inX <= "0000000000000000"; inY <= "1111111111111111";
      inZX <= '1'; inNX <= '1'; inZY <= '0'; inNY <= '0'; inF <= "00"; inNO <= '0'; inSizeX <= "000"; inSizeY <= "000"; inDirX <= '0'; inDirY <= '0';
      wait for 200 ps;
      assert(outZR = '0' and outNG = '1' and outSaida= "1111111111111111")  report "Falha em teste: 6" severity error;

      -- Teste: 7
      inX <= "0000000000000000"; inY <= "1111111111111111";
      inZX <= '0'; inNX <= '0'; inZY <= '1'; inNY <= '1'; inF <= "00"; inNO <= '1'; inSizeX <= "000"; inSizeY <= "000"; inDirX <= '0'; inDirY <= '0';
      wait for 200 ps;
      assert(outZR = '0' and outNG = '1' and outSaida= "1111111111111111")  report "Falha em teste: 7" severity error;

      -- Teste: 8
      inX <= "0000000000000000"; inY <= "1111111111111111";
      inZX <= '1'; inNX <= '1'; inZY <= '0'; inNY <= '0'; inF <= "00"; inNO <= '1'; inSizeX <= "000"; inSizeY <= "000"; inDirX <= '0'; inDirY <= '0';
      wait for 200 ps;
      assert(outZR = '1' and outNG = '0' and outSaida= "0000000000000000")  report "Falha em teste: 8" severity error;

      -- Teste: 9
      inX <= "0000000000000000"; inY <= "1111111111111111";
      inZX <= '0'; inNX <= '0'; inZY <= '1'; inNY <= '1'; inF <= "01"; inNO <= '1'; inSizeX <= "000"; inSizeY <= "000"; inDirX <= '0'; inDirY <= '0';
      wait for 200 ps;
      assert(outZR = '1' and outNG = '0' and outSaida= "0000000000000000")  report "Falha em teste: 9" severity error;

      -- Teste: 10
      inX <= "0000000000000000"; inY <= "1111111111111111";
      inZX <= '1'; inNX <= '1'; inZY <= '0'; inNY <= '0'; inF <= "01"; inNO <= '1'; inSizeX <= "000"; inSizeY <= "000"; inDirX <= '0'; inDirY <= '0';
      wait for 200 ps;
      assert(outZR = '0' and outNG = '0' and outSaida= "0000000000000001")  report "Falha em teste: 10" severity error;

      -- Teste: 11
      inX <= "0000000000000000"; inY <= "1111111111111111";
      inZX <= '0'; inNX <= '1'; inZY <= '1'; inNY <= '1'; inF <= "01"; inNO <= '1'; inSizeX <= "000"; inSizeY <= "000"; inDirX <= '0'; inDirY <= '0';
      wait for 200 ps;
      assert(outZR = '0' and outNG = '0' and outSaida= "0000000000000001")  report "Falha em teste: 11" severity error;

      -- Teste: 12
      inX <= "0000000000000000"; inY <= "1111111111111111";
      inZX <= '1'; inNX <= '1'; inZY <= '0'; inNY <= '1'; inF <= "01"; inNO <= '1'; inSizeX <= "000"; inSizeY <= "000"; inDirX <= '0'; inDirY <= '0';
      wait for 200 ps;
      assert(outZR = '1' and outNG = '0' and outSaida= "0000000000000000")  report "Falha em teste: 12" severity error;

      -- Teste: 13
      inX <= "0000000000000000"; inY <= "1111111111111111";
      inZX <= '0'; inNX <= '0'; inZY <= '1'; inNY <= '1'; inF <= "01"; inNO <= '0'; inSizeX <= "000"; inSizeY <= "000"; inDirX <= '0'; inDirY <= '0';
      wait for 200 ps;
      assert(outZR = '0' and outNG = '1' and outSaida= "1111111111111111")  report "Falha em teste: 13" severity error;

      -- Teste: 14
      inX <= "0000000000000000"; inY <= "1111111111111111";
      inZX <= '1'; inNX <= '1'; inZY <= '0'; inNY <= '0'; inF <= "01"; inNO <= '0'; inSizeX <= "000"; inSizeY <= "000"; inDirX <= '0'; inDirY <= '0';
      wait for 200 ps;
      assert(outZR = '0' and outNG = '1' and outSaida= "1111111111111110")  report "Falha em teste: 14" severity error;

      -- Teste: 15
      inX <= "0000000000000000"; inY <= "1111111111111111";
      inZX <= '0'; inNX <= '0'; inZY <= '0'; inNY <= '0'; inF <= "01"; inNO <= '0'; inSizeX <= "000"; inSizeY <= "000"; inDirX <= '0'; inDirY <= '0';
      wait for 200 ps;
      assert(outZR = '0' and outNG = '1' and outSaida= "1111111111111111")  report "Falha em teste: 15" severity error;

      -- Teste: 16
      inX <= "0000000000000000"; inY <= "1111111111111111";
      inZX <= '0'; inNX <= '1'; inZY <= '0'; inNY <= '0'; inF <= "01"; inNO <= '1'; inSizeX <= "000"; inSizeY <= "000"; inDirX <= '0'; inDirY <= '0';
      wait for 200 ps;
      assert(outZR = '0' and outNG = '0' and outSaida= "0000000000000001")  report "Falha em teste: 16" severity error;

      -- Teste: 17
      inX <= "0000000000000000"; inY <= "1111111111111111";
      inZX <= '0'; inNX <= '0'; inZY <= '0'; inNY <= '1'; inF <= "01"; inNO <= '1'; inSizeX <= "000"; inSizeY <= "000"; inDirX <= '0'; inDirY <= '0';
      wait for 200 ps;
      assert(outZR = '0' and outNG = '1' and outSaida= "1111111111111111")  report "Falha em teste: 17" severity error;

      -- Teste: 18
      inX <= "0000000000000000"; inY <= "1111111111111111";
      inZX <= '0'; inNX <= '0'; inZY <= '0'; inNY <= '0'; inF <= "00"; inNO <= '0'; inSizeX <= "000"; inSizeY <= "000"; inDirX <= '0'; inDirY <= '0';
      wait for 200 ps;
      assert(outZR = '1' and outNG = '0' and outSaida= "0000000000000000")  report "Falha em teste: 18" severity error;

      -- Teste: 19
      inX <= "0000000000000000"; inY <= "1111111111111111";
      inZX <= '0'; inNX <= '1'; inZY <= '0'; inNY <= '1'; inF <= "00"; inNO <= '1'; inSizeX <= "000"; inSizeY <= "000"; inDirX <= '0'; inDirY <= '0';
      wait for 200 ps;
      assert(outZR = '0' and outNG = '1' and outSaida= "1111111111111111")  report "Falha em teste: 19" severity error;

      -- Teste: 20 (XOR)
      inX <= "0000000000000000"; inY <= "1111111111111111";
      inZX <= '0'; inNX <= '0'; inZY <= '0'; inNY <= '0'; inF <= "10"; inNO <= '0'; inSizeX <= "000"; inSizeY <= "000"; inDirX <= '0'; inDirY <= '0';
      wait for 200 ps;
      assert(outZR = '0' and outNG = '1' and outSaida= "1111111111111111")  report "Falha em teste: 20 (XOR)" severity error;

      -- Teste: 21 (XOR)
      inX <= "0011100100111000"; inY <= "0110101100101000";
      inZX <= '0'; inNX <= '0'; inZY <= '0'; inNY <= '0'; inF <= "10"; inNO <= '0'; inSizeX <= "000"; inSizeY <= "000"; inDirX <= '0'; inDirY <= '0';
      wait for 200 ps;
      assert(outZR = '0' and outNG = '0' and outSaida= "0101001000010000")  report "Falha em teste: 21 (XOR)" severity error;

      -- Teste: 22 (CARRY)
      inX <= "0000000000000001"; inY <= "1111111111111111";
      inZX <= '0'; inNX <= '0'; inZY <= '0'; inNY <= '0'; inF <= "01"; inNO <= '0'; inSizeX <= "000"; inSizeY <= "000"; inDirX <= '0'; inDirY <= '0';
      wait for 200 ps;
      assert(outZR = '1' and outNG = '0' and outSaida= "0000000000000000" and outCa='1')  report "Falha em teste: 22 (XOR)" severity error;

      -- Teste: 23 (CARRY)
      inX <= "0000000000000001"; inY <= "0000000000000001";
      inZX <= '0'; inNX <= '0'; inZY <= '0'; inNY <= '0'; inF <= "01"; inNO <= '0'; inSizeX <= "000"; inSizeY <= "000"; inDirX <= '0'; inDirY <= '0';
      wait for 200 ps;
      assert(outZR = '0' and outNG = '0' and outSaida= "0000000000000010" and outCa='0')  report "Falha em teste: 23 (XOR)" severity error;

      -- Teste: 24 (SHIFTER RIGHT)
      inX <= "0100000000000000"; inY <= "0100000000000000";
      inZX <= '0'; inNX <= '0'; inZY <= '0'; inNY <= '0'; inF <= "01"; inNO <= '0'; inSizeX <= "011"; inSizeY <= "100"; inDirX <= '1'; inDirY <= '1';
      wait for 200 ps;
      assert(outZR = '0' and outNG = '0' and outSaida= "0000110000000000" and outCa='0')  report "Falha em teste: Teste: 24 (SHIFTER RIGHT)" severity error;

      -- Teste: 23 (SHIFTER LEFT)
      inX <= "0000000000000010"; inY <= "0000000000000010";
      inZX <= '0'; inNX <= '0'; inZY <= '0'; inNY <= '0'; inF <= "01"; inNO <= '0'; inSizeX <= "000"; inSizeY <= "001"; inDirX <= '0'; inDirY <= '0';
      wait for 200 ps;
      assert(outZR = '0' and outNG = '0' and outSaida= "0000000000000110" and outCa='0')  report "Falha em teste: 23 (SHIFTER LEFT)" severity error;

    test_runner_cleanup(runner); -- Simulacao acaba aqui

  end process;
end architecture;
